package top_pkg;
		`include "uvm_macros.svh"

		import uvm_pkg::* ;
		import apb_pkg::* ;

		`include "scoreboard.sv"
		`include "environment_config.sv"
		`include "environment.sv"
		`include "base_test.sv"
		`include "sequence_library.sv"
		`include "test_library.sv"



endpackage


