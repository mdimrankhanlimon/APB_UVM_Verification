`include "reset_seq.sv"
`include "error_drive_seq.sv"
`include "cont_wr_rd_seq.sv"
`include "sanity_simple_seq.sv"

`include "cont_wr_rd_knobs_seq.sv"

`include "c_wr_rd_byte_ALinc_seq.sv"
`include "cont_wr_rd_knobs_loc_seq.sv"
