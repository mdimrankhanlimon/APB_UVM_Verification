`define    DEPTH 1024 
`define    ADDR_WIDTH $clog2(`DEPTH)
`define    DATA_WIDTH 32
`define    BYTE_LANE 4
