`include "apb_interface.sv"


package apb_pkg;
		`include "uvm_macros.svh"

		import uvm_pkg::* ;


		`include "apb_defines.sv"
		`include "apb_seq_item.sv"
		`include "apb_seq_lib.sv"
		`include "apb_sequencer.sv"
		`include "apb_driver_callback.sv"
		`include "apb_driver.sv"
		`include "apb_monitor.sv"
		`include "apb_coverage.sv"
		`include "apb_agent_config.sv"
		`include "apb_agent.sv"



endpackage

