//`include "base_test.sv"
`include "sanity_simple_test.sv"
`include "cont_wr_rd_test.sv"

`include "c_wr_rd_knobs_loc_test.sv"

`include "error_test.sv"
`include "reset_test.sv"

`include "c_wr_rd_byte_test.sv"
